`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory  
// Module - PCAdder.v
// Description - 32-Bit program counter (PC) adder.
// 
// INPUTS:-
// PCResult: 32-Bit input port.
// 
// OUTPUTS:-
// PCAddResult: 32-Bit output port.
//
// FUNCTIONALITY:-
// Design an incrementor (or a hard-wired ADD ALU whose first input is from the 
// PC, and whose second input is a hard-wired 4) that computes the current 
// PC + 4. The result should always be an increment of the signal 'PCResult' by 
// 4 (i.e., PCAddResult = PCResult + 4).
////////////////////////////////////////////////////////////////////////////////

module ProgramCounter(PCIn, PCOut,Clk,Reset,PCWrite);

    input [31:0] PCIn;
    input Clk;
    input Reset;
    input PCWrite;
   
    
    
    output reg [31:0] PCOut;
   
      
    
    
    always @(posedge Clk or posedge Reset) begin
        if ( Reset == 1) begin

                PCOut <= 0;
            end
        
            else if (PCWrite != 1)  begin
                PCOut <= PCIn;
            end
       
    end
    
endmodule

